// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II 64-Bit"
// VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"
// CREATED		"Mon May 02 20:12:52 2022"

module EXP33(
	CLK,
	ax_v,
	cx_v,
	IMM_v,
	MAR_v,
	PC_v,
	upc
);


input wire	CLK;
output wire	[15:0] ax_v;
output wire	[15:0] cx_v;
output wire	[15:0] IMM_v;
output wire	[7:0] MAR_v;
output wire	[15:0] PC_v;
output wire	[7:0] upc;

wire	[5:0] ALUOP;
wire	[15:0] BUSLINE;
wire	DBG1;
wire	DBG2;
wire	DBG3;
wire	DBG4;
wire	DBG5;
wire	DBG6;
wire	halo;
wire	[15:0] irb;
wire	[15:0] MARB;
wire	RDPC;
wire	[15:0] SPAB;
wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_62;
wire	SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_7;
wire	[2:0] SYNTHESIZED_WIRE_63;
wire	[2:0] SYNTHESIZED_WIRE_64;
wire	[2:0] SYNTHESIZED_WIRE_65;
wire	[3:0] SYNTHESIZED_WIRE_12;
wire	[3:0] SYNTHESIZED_WIRE_16;
wire	SYNTHESIZED_WIRE_17;
wire	SYNTHESIZED_WIRE_18;
wire	SYNTHESIZED_WIRE_20;
wire	SYNTHESIZED_WIRE_66;
wire	[7:0] SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_24;
wire	SYNTHESIZED_WIRE_25;
reg	DFF_odff;
wire	SYNTHESIZED_WIRE_26;
wire	SYNTHESIZED_WIRE_27;
wire	[2:0] SYNTHESIZED_WIRE_28;
wire	[15:0] SYNTHESIZED_WIRE_29;
wire	[15:0] SYNTHESIZED_WIRE_30;
wire	[15:0] SYNTHESIZED_WIRE_31;
wire	SYNTHESIZED_WIRE_32;
wire	[15:0] SYNTHESIZED_WIRE_33;
wire	SYNTHESIZED_WIRE_34;
wire	[15:0] SYNTHESIZED_WIRE_35;
wire	SYNTHESIZED_WIRE_36;
wire	SYNTHESIZED_WIRE_37;
wire	SYNTHESIZED_WIRE_38;
wire	SYNTHESIZED_WIRE_40;
wire	SYNTHESIZED_WIRE_42;
wire	SYNTHESIZED_WIRE_44;
wire	SYNTHESIZED_WIRE_45;
wire	SYNTHESIZED_WIRE_47;
wire	SYNTHESIZED_WIRE_48;
wire	SYNTHESIZED_WIRE_50;
wire	SYNTHESIZED_WIRE_51;
wire	SYNTHESIZED_WIRE_53;
wire	SYNTHESIZED_WIRE_54;
wire	SYNTHESIZED_WIRE_56;
wire	SYNTHESIZED_WIRE_57;
wire	SYNTHESIZED_WIRE_59;
wire	SYNTHESIZED_WIRE_60;

assign	SYNTHESIZED_WIRE_38 = 0;
assign	SYNTHESIZED_WIRE_40 = 1;
assign	SYNTHESIZED_WIRE_45 = 1;
assign	SYNTHESIZED_WIRE_51 = 0;




REG16-TRI-IMM-BN	b2v_BX(
	.WN(SYNTHESIZED_WIRE_0),
	.RN(SYNTHESIZED_WIRE_1),
	.CLK(SYNTHESIZED_WIRE_62),
	.D(BUSLINE),
	
	.Otri(BUSLINE));


REG16-TRI-IMM-BN	b2v_CX(
	.WN(SYNTHESIZED_WIRE_3),
	.RN(SYNTHESIZED_WIRE_4),
	.CLK(SYNTHESIZED_WIRE_62),
	.D(BUSLINE),
	.Oimm(cx_v),
	.Otri(BUSLINE));


REG16-TRI-IMM-BN	b2v_DX(
	.WN(SYNTHESIZED_WIRE_6),
	.RN(SYNTHESIZED_WIRE_7),
	.CLK(SYNTHESIZED_WIRE_62),
	.D(BUSLINE),
	
	.Otri(BUSLINE));


FINDER	b2v_FINDER-READ(
	.R1(SYNTHESIZED_WIRE_63),
	.R2(SYNTHESIZED_WIRE_64),
	.R3(SYNTHESIZED_WIRE_65),
	.SY(SYNTHESIZED_WIRE_12),
	.AXN(SYNTHESIZED_WIRE_48),
	.BXN(SYNTHESIZED_WIRE_1),
	.CXN(SYNTHESIZED_WIRE_4),
	.DXN(SYNTHESIZED_WIRE_7),
	.SPAN(SYNTHESIZED_WIRE_54),
	.SPBN(SYNTHESIZED_WIRE_57),
	.SPCN(SYNTHESIZED_WIRE_60),
	.IMMN(SYNTHESIZED_WIRE_18),
	.PCN(RDPC),
	
	
	
	.alu_lN(SYNTHESIZED_WIRE_27),
	.alu_hN(SYNTHESIZED_WIRE_26),
	.RAMN(SYNTHESIZED_WIRE_24));


FINDER	b2v_FINDER-WRITE(
	.R1(SYNTHESIZED_WIRE_63),
	.R2(SYNTHESIZED_WIRE_64),
	.R3(SYNTHESIZED_WIRE_65),
	.SY(SYNTHESIZED_WIRE_16),
	.AXN(SYNTHESIZED_WIRE_47),
	.BXN(SYNTHESIZED_WIRE_0),
	.CXN(SYNTHESIZED_WIRE_3),
	.DXN(SYNTHESIZED_WIRE_6),
	.SPAN(SYNTHESIZED_WIRE_53),
	.SPBN(SYNTHESIZED_WIRE_56),
	.SPCN(SYNTHESIZED_WIRE_59),
	.IMMN(SYNTHESIZED_WIRE_17),
	.PCN(SYNTHESIZED_WIRE_42),
	.MARN(SYNTHESIZED_WIRE_37),
	
	.IRN(SYNTHESIZED_WIRE_50),
	
	
	.RAMN(SYNTHESIZED_WIRE_25));


REG16-TRI-IMM-BN	b2v_imm(
	.WN(SYNTHESIZED_WIRE_17),
	.RN(SYNTHESIZED_WIRE_18),
	.CLK(SYNTHESIZED_WIRE_62),
	.D(BUSLINE),
	.Oimm(IMM_v),
	.Otri(BUSLINE));


CU	b2v_inst(
	.immE(SYNTHESIZED_WIRE_20),
	.CLK(SYNTHESIZED_WIRE_66),
	.iAddr(SYNTHESIZED_WIRE_22),
	.halt(halo),
	.ALU_ENA(SYNTHESIZED_WIRE_28),
	.ALU_OP(ALUOP),
	.DBG_UPC(upc),
	.READ(SYNTHESIZED_WIRE_12),
	.WRITE(SYNTHESIZED_WIRE_16));

assign	SYNTHESIZED_WIRE_62 =  ~SYNTHESIZED_WIRE_66;

assign	SYNTHESIZED_WIRE_36 =  ~SYNTHESIZED_WIRE_24;

assign	SYNTHESIZED_WIRE_44 =  ~SYNTHESIZED_WIRE_25;

assign	SYNTHESIZED_WIRE_66 = CLK | DFF_odff;



assign	SYNTHESIZED_WIRE_34 =  ~SYNTHESIZED_WIRE_26;


assign	SYNTHESIZED_WIRE_32 =  ~SYNTHESIZED_WIRE_27;


ALU16	b2v_inst4(
	.ENA(SYNTHESIZED_WIRE_28),
	.OP(ALUOP),
	.SPA(SPAB),
	.SPB(SYNTHESIZED_WIRE_29),
	.SPC(SYNTHESIZED_WIRE_30),
	
	
	
	
	
	
	.OUTH(SYNTHESIZED_WIRE_33),
	.OUTL(SYNTHESIZED_WIRE_31));


assign	BUSLINE[15] = SYNTHESIZED_WIRE_32 ? SYNTHESIZED_WIRE_31[15] : 1'bz;
assign	BUSLINE[14] = SYNTHESIZED_WIRE_32 ? SYNTHESIZED_WIRE_31[14] : 1'bz;
assign	BUSLINE[13] = SYNTHESIZED_WIRE_32 ? SYNTHESIZED_WIRE_31[13] : 1'bz;
assign	BUSLINE[12] = SYNTHESIZED_WIRE_32 ? SYNTHESIZED_WIRE_31[12] : 1'bz;
assign	BUSLINE[11] = SYNTHESIZED_WIRE_32 ? SYNTHESIZED_WIRE_31[11] : 1'bz;
assign	BUSLINE[10] = SYNTHESIZED_WIRE_32 ? SYNTHESIZED_WIRE_31[10] : 1'bz;
assign	BUSLINE[9] = SYNTHESIZED_WIRE_32 ? SYNTHESIZED_WIRE_31[9] : 1'bz;
assign	BUSLINE[8] = SYNTHESIZED_WIRE_32 ? SYNTHESIZED_WIRE_31[8] : 1'bz;
assign	BUSLINE[7] = SYNTHESIZED_WIRE_32 ? SYNTHESIZED_WIRE_31[7] : 1'bz;
assign	BUSLINE[6] = SYNTHESIZED_WIRE_32 ? SYNTHESIZED_WIRE_31[6] : 1'bz;
assign	BUSLINE[5] = SYNTHESIZED_WIRE_32 ? SYNTHESIZED_WIRE_31[5] : 1'bz;
assign	BUSLINE[4] = SYNTHESIZED_WIRE_32 ? SYNTHESIZED_WIRE_31[4] : 1'bz;
assign	BUSLINE[3] = SYNTHESIZED_WIRE_32 ? SYNTHESIZED_WIRE_31[3] : 1'bz;
assign	BUSLINE[2] = SYNTHESIZED_WIRE_32 ? SYNTHESIZED_WIRE_31[2] : 1'bz;
assign	BUSLINE[1] = SYNTHESIZED_WIRE_32 ? SYNTHESIZED_WIRE_31[1] : 1'bz;
assign	BUSLINE[0] = SYNTHESIZED_WIRE_32 ? SYNTHESIZED_WIRE_31[0] : 1'bz;

assign	BUSLINE[15] = SYNTHESIZED_WIRE_34 ? SYNTHESIZED_WIRE_33[15] : 1'bz;
assign	BUSLINE[14] = SYNTHESIZED_WIRE_34 ? SYNTHESIZED_WIRE_33[14] : 1'bz;
assign	BUSLINE[13] = SYNTHESIZED_WIRE_34 ? SYNTHESIZED_WIRE_33[13] : 1'bz;
assign	BUSLINE[12] = SYNTHESIZED_WIRE_34 ? SYNTHESIZED_WIRE_33[12] : 1'bz;
assign	BUSLINE[11] = SYNTHESIZED_WIRE_34 ? SYNTHESIZED_WIRE_33[11] : 1'bz;
assign	BUSLINE[10] = SYNTHESIZED_WIRE_34 ? SYNTHESIZED_WIRE_33[10] : 1'bz;
assign	BUSLINE[9] = SYNTHESIZED_WIRE_34 ? SYNTHESIZED_WIRE_33[9] : 1'bz;
assign	BUSLINE[8] = SYNTHESIZED_WIRE_34 ? SYNTHESIZED_WIRE_33[8] : 1'bz;
assign	BUSLINE[7] = SYNTHESIZED_WIRE_34 ? SYNTHESIZED_WIRE_33[7] : 1'bz;
assign	BUSLINE[6] = SYNTHESIZED_WIRE_34 ? SYNTHESIZED_WIRE_33[6] : 1'bz;
assign	BUSLINE[5] = SYNTHESIZED_WIRE_34 ? SYNTHESIZED_WIRE_33[5] : 1'bz;
assign	BUSLINE[4] = SYNTHESIZED_WIRE_34 ? SYNTHESIZED_WIRE_33[4] : 1'bz;
assign	BUSLINE[3] = SYNTHESIZED_WIRE_34 ? SYNTHESIZED_WIRE_33[3] : 1'bz;
assign	BUSLINE[2] = SYNTHESIZED_WIRE_34 ? SYNTHESIZED_WIRE_33[2] : 1'bz;
assign	BUSLINE[1] = SYNTHESIZED_WIRE_34 ? SYNTHESIZED_WIRE_33[1] : 1'bz;
assign	BUSLINE[0] = SYNTHESIZED_WIRE_34 ? SYNTHESIZED_WIRE_33[0] : 1'bz;


DECODER	b2v_inst8(
	.IR(irb),
	.immE(SYNTHESIZED_WIRE_20),
	.R1(SYNTHESIZED_WIRE_63),
	.R2(SYNTHESIZED_WIRE_64),
	.R3(SYNTHESIZED_WIRE_65),
	.uaddr(SYNTHESIZED_WIRE_22));

assign	BUSLINE[15] = SYNTHESIZED_WIRE_36 ? SYNTHESIZED_WIRE_35[15] : 1'bz;
assign	BUSLINE[14] = SYNTHESIZED_WIRE_36 ? SYNTHESIZED_WIRE_35[14] : 1'bz;
assign	BUSLINE[13] = SYNTHESIZED_WIRE_36 ? SYNTHESIZED_WIRE_35[13] : 1'bz;
assign	BUSLINE[12] = SYNTHESIZED_WIRE_36 ? SYNTHESIZED_WIRE_35[12] : 1'bz;
assign	BUSLINE[11] = SYNTHESIZED_WIRE_36 ? SYNTHESIZED_WIRE_35[11] : 1'bz;
assign	BUSLINE[10] = SYNTHESIZED_WIRE_36 ? SYNTHESIZED_WIRE_35[10] : 1'bz;
assign	BUSLINE[9] = SYNTHESIZED_WIRE_36 ? SYNTHESIZED_WIRE_35[9] : 1'bz;
assign	BUSLINE[8] = SYNTHESIZED_WIRE_36 ? SYNTHESIZED_WIRE_35[8] : 1'bz;
assign	BUSLINE[7] = SYNTHESIZED_WIRE_36 ? SYNTHESIZED_WIRE_35[7] : 1'bz;
assign	BUSLINE[6] = SYNTHESIZED_WIRE_36 ? SYNTHESIZED_WIRE_35[6] : 1'bz;
assign	BUSLINE[5] = SYNTHESIZED_WIRE_36 ? SYNTHESIZED_WIRE_35[5] : 1'bz;
assign	BUSLINE[4] = SYNTHESIZED_WIRE_36 ? SYNTHESIZED_WIRE_35[4] : 1'bz;
assign	BUSLINE[3] = SYNTHESIZED_WIRE_36 ? SYNTHESIZED_WIRE_35[3] : 1'bz;
assign	BUSLINE[2] = SYNTHESIZED_WIRE_36 ? SYNTHESIZED_WIRE_35[2] : 1'bz;
assign	BUSLINE[1] = SYNTHESIZED_WIRE_36 ? SYNTHESIZED_WIRE_35[1] : 1'bz;
assign	BUSLINE[0] = SYNTHESIZED_WIRE_36 ? SYNTHESIZED_WIRE_35[0] : 1'bz;


REG16-TRI-B-N	b2v_MAR(
	.WN(SYNTHESIZED_WIRE_37),
	.RN(SYNTHESIZED_WIRE_38),
	.CLK(SYNTHESIZED_WIRE_62),
	.I(BUSLINE),
	.O(MARB));


always@(posedge SYNTHESIZED_WIRE_62 or negedge SYNTHESIZED_WIRE_40)
begin
if (!SYNTHESIZED_WIRE_40)
	begin
	DFF_odff <= 0;
	end
else
	begin
	DFF_odff <= halo;
	end
end


REG16-TRI-IMM-BN	b2v_PC(
	.WN(SYNTHESIZED_WIRE_42),
	.RN(RDPC),
	.CLK(SYNTHESIZED_WIRE_62),
	.D(BUSLINE),
	.Oimm(PC_v),
	.Otri(BUSLINE));


RAM0	b2v_RAM(
	.wren(SYNTHESIZED_WIRE_44),
	.rden(SYNTHESIZED_WIRE_45),
	.inclock(SYNTHESIZED_WIRE_62),
	.address(MARB[7:0]),
	.data(BUSLINE),
	.q(SYNTHESIZED_WIRE_35));


REG16-TRI-IMM-BN	b2v_reg-ax(
	.WN(SYNTHESIZED_WIRE_47),
	.RN(SYNTHESIZED_WIRE_48),
	.CLK(SYNTHESIZED_WIRE_62),
	.D(BUSLINE),
	.Oimm(ax_v),
	.Otri(BUSLINE));


REG16-TRI-B-N	b2v_reg-ir(
	.WN(SYNTHESIZED_WIRE_50),
	.RN(SYNTHESIZED_WIRE_51),
	.CLK(SYNTHESIZED_WIRE_62),
	.I(BUSLINE),
	.O(irb));


REG16-TRI-IMM-BN	b2v_spA(
	.WN(SYNTHESIZED_WIRE_53),
	.RN(SYNTHESIZED_WIRE_54),
	.CLK(SYNTHESIZED_WIRE_62),
	.D(BUSLINE),
	.Oimm(SPAB),
	.Otri(BUSLINE));


REG16-TRI-IMM-BN	b2v_spB(
	.WN(SYNTHESIZED_WIRE_56),
	.RN(SYNTHESIZED_WIRE_57),
	.CLK(SYNTHESIZED_WIRE_62),
	.D(BUSLINE),
	.Oimm(SYNTHESIZED_WIRE_29),
	.Otri(BUSLINE));


REG16-TRI-IMM-BN	b2v_spC(
	.WN(SYNTHESIZED_WIRE_59),
	.RN(SYNTHESIZED_WIRE_60),
	.CLK(SYNTHESIZED_WIRE_62),
	.D(BUSLINE),
	.Oimm(SYNTHESIZED_WIRE_30),
	.Otri(BUSLINE));

assign	MAR_v[7:0] = MARB[7:0];

endmodule
