-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"
-- CREATED		"Mon May 02 20:12:02 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY EXP33 IS 
	PORT
	(
		CLK :  IN  STD_LOGIC;
		ax_v :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		cx_v :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		IMM_v :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		MAR_v :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		PC_v :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		upc :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END EXP33;

ARCHITECTURE bdf_type OF EXP33 IS 

COMPONENT reg16-tri-imm-bn
	PORT(WN : IN STD_LOGIC;
		 RN : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 D : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 Oimm : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 Otri : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT finder
	PORT(R1 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 R2 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 R3 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 SY : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 AXN : OUT STD_LOGIC;
		 BXN : OUT STD_LOGIC;
		 CXN : OUT STD_LOGIC;
		 DXN : OUT STD_LOGIC;
		 SPAN : OUT STD_LOGIC;
		 SPBN : OUT STD_LOGIC;
		 SPCN : OUT STD_LOGIC;
		 IMMN : OUT STD_LOGIC;
		 PCN : OUT STD_LOGIC;
		 MARN : OUT STD_LOGIC;
		 MDRN : OUT STD_LOGIC;
		 IRN : OUT STD_LOGIC;
		 alu_lN : OUT STD_LOGIC;
		 alu_hN : OUT STD_LOGIC;
		 RAMN : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT cu
	PORT(immE : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 iAddr : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 halt : OUT STD_LOGIC;
		 ALU_ENA : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		 ALU_OP : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		 DBG_UPC : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 READ : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 WRITE : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT alu16
	PORT(ENA : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 OP : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 SPA : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 SPB : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 SPC : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 DBG1 : OUT STD_LOGIC;
		 DBG2 : OUT STD_LOGIC;
		 DBG3 : OUT STD_LOGIC;
		 DBG4 : OUT STD_LOGIC;
		 DBG5 : OUT STD_LOGIC;
		 DBG6 : OUT STD_LOGIC;
		 OUTH : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 OUTL : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT decoder
	PORT(IR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 immE : OUT STD_LOGIC;
		 R1 : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		 R2 : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		 R3 : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		 uaddr : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT reg16-tri-b-n
	PORT(WN : IN STD_LOGIC;
		 RN : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 I : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 O : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ram0
	PORT(wren : IN STD_LOGIC;
		 rden : IN STD_LOGIC;
		 inclock : IN STD_LOGIC;
		 address : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 data : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	ALUOP :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	BUSLINE :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	DBG1 :  STD_LOGIC;
SIGNAL	DBG2 :  STD_LOGIC;
SIGNAL	DBG3 :  STD_LOGIC;
SIGNAL	DBG4 :  STD_LOGIC;
SIGNAL	DBG5 :  STD_LOGIC;
SIGNAL	DBG6 :  STD_LOGIC;
SIGNAL	halo :  STD_LOGIC;
SIGNAL	irb :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	MARB :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	RDPC :  STD_LOGIC;
SIGNAL	SPAB :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	DFF_odff :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_41 <= '0';
SYNTHESIZED_WIRE_44 <= '0';
SYNTHESIZED_WIRE_46 <= '1';
SYNTHESIZED_WIRE_51 <= '1';



b2v_AX : reg16-tri-imm-bn
PORT MAP(WN => SYNTHESIZED_WIRE_0,
		 RN => SYNTHESIZED_WIRE_1,
		 CLK => SYNTHESIZED_WIRE_62,
		 D => BUSLINE,
		 Oimm => ax_v,
		 Otri => BUSLINE);


b2v_BX : reg16-tri-imm-bn
PORT MAP(WN => SYNTHESIZED_WIRE_3,
		 RN => SYNTHESIZED_WIRE_4,
		 CLK => SYNTHESIZED_WIRE_62,
		 D => BUSLINE,
		 Otri => BUSLINE);


b2v_CX : reg16-tri-imm-bn
PORT MAP(WN => SYNTHESIZED_WIRE_6,
		 RN => SYNTHESIZED_WIRE_7,
		 CLK => SYNTHESIZED_WIRE_62,
		 D => BUSLINE,
		 Oimm => cx_v,
		 Otri => BUSLINE);


b2v_DX : reg16-tri-imm-bn
PORT MAP(WN => SYNTHESIZED_WIRE_9,
		 RN => SYNTHESIZED_WIRE_10,
		 CLK => SYNTHESIZED_WIRE_62,
		 D => BUSLINE,
		 Otri => BUSLINE);


b2v_FINDER-READ : finder
PORT MAP(R1 => SYNTHESIZED_WIRE_63,
		 R2 => SYNTHESIZED_WIRE_64,
		 R3 => SYNTHESIZED_WIRE_65,
		 SY => SYNTHESIZED_WIRE_15,
		 AXN => SYNTHESIZED_WIRE_1,
		 BXN => SYNTHESIZED_WIRE_4,
		 CXN => SYNTHESIZED_WIRE_7,
		 DXN => SYNTHESIZED_WIRE_10,
		 SPAN => SYNTHESIZED_WIRE_54,
		 SPBN => SYNTHESIZED_WIRE_57,
		 SPCN => SYNTHESIZED_WIRE_60,
		 IMMN => SYNTHESIZED_WIRE_21,
		 PCN => RDPC,
		 alu_lN => SYNTHESIZED_WIRE_30,
		 alu_hN => SYNTHESIZED_WIRE_29,
		 RAMN => SYNTHESIZED_WIRE_27);


b2v_FINDER-WRITE : finder
PORT MAP(R1 => SYNTHESIZED_WIRE_63,
		 R2 => SYNTHESIZED_WIRE_64,
		 R3 => SYNTHESIZED_WIRE_65,
		 SY => SYNTHESIZED_WIRE_19,
		 AXN => SYNTHESIZED_WIRE_0,
		 BXN => SYNTHESIZED_WIRE_3,
		 CXN => SYNTHESIZED_WIRE_6,
		 DXN => SYNTHESIZED_WIRE_9,
		 SPAN => SYNTHESIZED_WIRE_53,
		 SPBN => SYNTHESIZED_WIRE_56,
		 SPCN => SYNTHESIZED_WIRE_59,
		 IMMN => SYNTHESIZED_WIRE_20,
		 PCN => SYNTHESIZED_WIRE_48,
		 MARN => SYNTHESIZED_WIRE_43,
		 IRN => SYNTHESIZED_WIRE_40,
		 RAMN => SYNTHESIZED_WIRE_28);


b2v_imm : reg16-tri-imm-bn
PORT MAP(WN => SYNTHESIZED_WIRE_20,
		 RN => SYNTHESIZED_WIRE_21,
		 CLK => SYNTHESIZED_WIRE_62,
		 D => BUSLINE,
		 Oimm => IMM_v,
		 Otri => BUSLINE);


b2v_inst : cu
PORT MAP(immE => SYNTHESIZED_WIRE_23,
		 CLK => SYNTHESIZED_WIRE_66,
		 iAddr => SYNTHESIZED_WIRE_25,
		 halt => halo,
		 ALU_ENA => SYNTHESIZED_WIRE_31,
		 ALU_OP => ALUOP,
		 DBG_UPC => upc,
		 READ => SYNTHESIZED_WIRE_15,
		 WRITE => SYNTHESIZED_WIRE_19);


SYNTHESIZED_WIRE_62 <= NOT(SYNTHESIZED_WIRE_66);



SYNTHESIZED_WIRE_39 <= NOT(SYNTHESIZED_WIRE_27);



SYNTHESIZED_WIRE_50 <= NOT(SYNTHESIZED_WIRE_28);



SYNTHESIZED_WIRE_66 <= CLK OR DFF_odff;




SYNTHESIZED_WIRE_37 <= NOT(SYNTHESIZED_WIRE_29);




SYNTHESIZED_WIRE_35 <= NOT(SYNTHESIZED_WIRE_30);



b2v_inst4 : alu16
PORT MAP(ENA => SYNTHESIZED_WIRE_31,
		 OP => ALUOP,
		 SPA => SPAB,
		 SPB => SYNTHESIZED_WIRE_32,
		 SPC => SYNTHESIZED_WIRE_33,
		 OUTH => SYNTHESIZED_WIRE_36,
		 OUTL => SYNTHESIZED_WIRE_34);



PROCESS(SYNTHESIZED_WIRE_34,SYNTHESIZED_WIRE_35)
BEGIN
if (SYNTHESIZED_WIRE_35 = '1') THEN
	BUSLINE(15) <= SYNTHESIZED_WIRE_34(15);
ELSE
	BUSLINE(15) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_34,SYNTHESIZED_WIRE_35)
BEGIN
if (SYNTHESIZED_WIRE_35 = '1') THEN
	BUSLINE(14) <= SYNTHESIZED_WIRE_34(14);
ELSE
	BUSLINE(14) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_34,SYNTHESIZED_WIRE_35)
BEGIN
if (SYNTHESIZED_WIRE_35 = '1') THEN
	BUSLINE(13) <= SYNTHESIZED_WIRE_34(13);
ELSE
	BUSLINE(13) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_34,SYNTHESIZED_WIRE_35)
BEGIN
if (SYNTHESIZED_WIRE_35 = '1') THEN
	BUSLINE(12) <= SYNTHESIZED_WIRE_34(12);
ELSE
	BUSLINE(12) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_34,SYNTHESIZED_WIRE_35)
BEGIN
if (SYNTHESIZED_WIRE_35 = '1') THEN
	BUSLINE(11) <= SYNTHESIZED_WIRE_34(11);
ELSE
	BUSLINE(11) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_34,SYNTHESIZED_WIRE_35)
BEGIN
if (SYNTHESIZED_WIRE_35 = '1') THEN
	BUSLINE(10) <= SYNTHESIZED_WIRE_34(10);
ELSE
	BUSLINE(10) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_34,SYNTHESIZED_WIRE_35)
BEGIN
if (SYNTHESIZED_WIRE_35 = '1') THEN
	BUSLINE(9) <= SYNTHESIZED_WIRE_34(9);
ELSE
	BUSLINE(9) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_34,SYNTHESIZED_WIRE_35)
BEGIN
if (SYNTHESIZED_WIRE_35 = '1') THEN
	BUSLINE(8) <= SYNTHESIZED_WIRE_34(8);
ELSE
	BUSLINE(8) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_34,SYNTHESIZED_WIRE_35)
BEGIN
if (SYNTHESIZED_WIRE_35 = '1') THEN
	BUSLINE(7) <= SYNTHESIZED_WIRE_34(7);
ELSE
	BUSLINE(7) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_34,SYNTHESIZED_WIRE_35)
BEGIN
if (SYNTHESIZED_WIRE_35 = '1') THEN
	BUSLINE(6) <= SYNTHESIZED_WIRE_34(6);
ELSE
	BUSLINE(6) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_34,SYNTHESIZED_WIRE_35)
BEGIN
if (SYNTHESIZED_WIRE_35 = '1') THEN
	BUSLINE(5) <= SYNTHESIZED_WIRE_34(5);
ELSE
	BUSLINE(5) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_34,SYNTHESIZED_WIRE_35)
BEGIN
if (SYNTHESIZED_WIRE_35 = '1') THEN
	BUSLINE(4) <= SYNTHESIZED_WIRE_34(4);
ELSE
	BUSLINE(4) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_34,SYNTHESIZED_WIRE_35)
BEGIN
if (SYNTHESIZED_WIRE_35 = '1') THEN
	BUSLINE(3) <= SYNTHESIZED_WIRE_34(3);
ELSE
	BUSLINE(3) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_34,SYNTHESIZED_WIRE_35)
BEGIN
if (SYNTHESIZED_WIRE_35 = '1') THEN
	BUSLINE(2) <= SYNTHESIZED_WIRE_34(2);
ELSE
	BUSLINE(2) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_34,SYNTHESIZED_WIRE_35)
BEGIN
if (SYNTHESIZED_WIRE_35 = '1') THEN
	BUSLINE(1) <= SYNTHESIZED_WIRE_34(1);
ELSE
	BUSLINE(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_34,SYNTHESIZED_WIRE_35)
BEGIN
if (SYNTHESIZED_WIRE_35 = '1') THEN
	BUSLINE(0) <= SYNTHESIZED_WIRE_34(0);
ELSE
	BUSLINE(0) <= 'Z';
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_36,SYNTHESIZED_WIRE_37)
BEGIN
if (SYNTHESIZED_WIRE_37 = '1') THEN
	BUSLINE(15) <= SYNTHESIZED_WIRE_36(15);
ELSE
	BUSLINE(15) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_36,SYNTHESIZED_WIRE_37)
BEGIN
if (SYNTHESIZED_WIRE_37 = '1') THEN
	BUSLINE(14) <= SYNTHESIZED_WIRE_36(14);
ELSE
	BUSLINE(14) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_36,SYNTHESIZED_WIRE_37)
BEGIN
if (SYNTHESIZED_WIRE_37 = '1') THEN
	BUSLINE(13) <= SYNTHESIZED_WIRE_36(13);
ELSE
	BUSLINE(13) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_36,SYNTHESIZED_WIRE_37)
BEGIN
if (SYNTHESIZED_WIRE_37 = '1') THEN
	BUSLINE(12) <= SYNTHESIZED_WIRE_36(12);
ELSE
	BUSLINE(12) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_36,SYNTHESIZED_WIRE_37)
BEGIN
if (SYNTHESIZED_WIRE_37 = '1') THEN
	BUSLINE(11) <= SYNTHESIZED_WIRE_36(11);
ELSE
	BUSLINE(11) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_36,SYNTHESIZED_WIRE_37)
BEGIN
if (SYNTHESIZED_WIRE_37 = '1') THEN
	BUSLINE(10) <= SYNTHESIZED_WIRE_36(10);
ELSE
	BUSLINE(10) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_36,SYNTHESIZED_WIRE_37)
BEGIN
if (SYNTHESIZED_WIRE_37 = '1') THEN
	BUSLINE(9) <= SYNTHESIZED_WIRE_36(9);
ELSE
	BUSLINE(9) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_36,SYNTHESIZED_WIRE_37)
BEGIN
if (SYNTHESIZED_WIRE_37 = '1') THEN
	BUSLINE(8) <= SYNTHESIZED_WIRE_36(8);
ELSE
	BUSLINE(8) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_36,SYNTHESIZED_WIRE_37)
BEGIN
if (SYNTHESIZED_WIRE_37 = '1') THEN
	BUSLINE(7) <= SYNTHESIZED_WIRE_36(7);
ELSE
	BUSLINE(7) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_36,SYNTHESIZED_WIRE_37)
BEGIN
if (SYNTHESIZED_WIRE_37 = '1') THEN
	BUSLINE(6) <= SYNTHESIZED_WIRE_36(6);
ELSE
	BUSLINE(6) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_36,SYNTHESIZED_WIRE_37)
BEGIN
if (SYNTHESIZED_WIRE_37 = '1') THEN
	BUSLINE(5) <= SYNTHESIZED_WIRE_36(5);
ELSE
	BUSLINE(5) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_36,SYNTHESIZED_WIRE_37)
BEGIN
if (SYNTHESIZED_WIRE_37 = '1') THEN
	BUSLINE(4) <= SYNTHESIZED_WIRE_36(4);
ELSE
	BUSLINE(4) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_36,SYNTHESIZED_WIRE_37)
BEGIN
if (SYNTHESIZED_WIRE_37 = '1') THEN
	BUSLINE(3) <= SYNTHESIZED_WIRE_36(3);
ELSE
	BUSLINE(3) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_36,SYNTHESIZED_WIRE_37)
BEGIN
if (SYNTHESIZED_WIRE_37 = '1') THEN
	BUSLINE(2) <= SYNTHESIZED_WIRE_36(2);
ELSE
	BUSLINE(2) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_36,SYNTHESIZED_WIRE_37)
BEGIN
if (SYNTHESIZED_WIRE_37 = '1') THEN
	BUSLINE(1) <= SYNTHESIZED_WIRE_36(1);
ELSE
	BUSLINE(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_36,SYNTHESIZED_WIRE_37)
BEGIN
if (SYNTHESIZED_WIRE_37 = '1') THEN
	BUSLINE(0) <= SYNTHESIZED_WIRE_36(0);
ELSE
	BUSLINE(0) <= 'Z';
END IF;
END PROCESS;


b2v_inst8 : decoder
PORT MAP(IR => irb,
		 immE => SYNTHESIZED_WIRE_23,
		 R1 => SYNTHESIZED_WIRE_63,
		 R2 => SYNTHESIZED_WIRE_64,
		 R3 => SYNTHESIZED_WIRE_65,
		 uaddr => SYNTHESIZED_WIRE_25);


PROCESS(SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_39)
BEGIN
if (SYNTHESIZED_WIRE_39 = '1') THEN
	BUSLINE(15) <= SYNTHESIZED_WIRE_38(15);
ELSE
	BUSLINE(15) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_39)
BEGIN
if (SYNTHESIZED_WIRE_39 = '1') THEN
	BUSLINE(14) <= SYNTHESIZED_WIRE_38(14);
ELSE
	BUSLINE(14) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_39)
BEGIN
if (SYNTHESIZED_WIRE_39 = '1') THEN
	BUSLINE(13) <= SYNTHESIZED_WIRE_38(13);
ELSE
	BUSLINE(13) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_39)
BEGIN
if (SYNTHESIZED_WIRE_39 = '1') THEN
	BUSLINE(12) <= SYNTHESIZED_WIRE_38(12);
ELSE
	BUSLINE(12) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_39)
BEGIN
if (SYNTHESIZED_WIRE_39 = '1') THEN
	BUSLINE(11) <= SYNTHESIZED_WIRE_38(11);
ELSE
	BUSLINE(11) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_39)
BEGIN
if (SYNTHESIZED_WIRE_39 = '1') THEN
	BUSLINE(10) <= SYNTHESIZED_WIRE_38(10);
ELSE
	BUSLINE(10) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_39)
BEGIN
if (SYNTHESIZED_WIRE_39 = '1') THEN
	BUSLINE(9) <= SYNTHESIZED_WIRE_38(9);
ELSE
	BUSLINE(9) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_39)
BEGIN
if (SYNTHESIZED_WIRE_39 = '1') THEN
	BUSLINE(8) <= SYNTHESIZED_WIRE_38(8);
ELSE
	BUSLINE(8) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_39)
BEGIN
if (SYNTHESIZED_WIRE_39 = '1') THEN
	BUSLINE(7) <= SYNTHESIZED_WIRE_38(7);
ELSE
	BUSLINE(7) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_39)
BEGIN
if (SYNTHESIZED_WIRE_39 = '1') THEN
	BUSLINE(6) <= SYNTHESIZED_WIRE_38(6);
ELSE
	BUSLINE(6) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_39)
BEGIN
if (SYNTHESIZED_WIRE_39 = '1') THEN
	BUSLINE(5) <= SYNTHESIZED_WIRE_38(5);
ELSE
	BUSLINE(5) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_39)
BEGIN
if (SYNTHESIZED_WIRE_39 = '1') THEN
	BUSLINE(4) <= SYNTHESIZED_WIRE_38(4);
ELSE
	BUSLINE(4) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_39)
BEGIN
if (SYNTHESIZED_WIRE_39 = '1') THEN
	BUSLINE(3) <= SYNTHESIZED_WIRE_38(3);
ELSE
	BUSLINE(3) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_39)
BEGIN
if (SYNTHESIZED_WIRE_39 = '1') THEN
	BUSLINE(2) <= SYNTHESIZED_WIRE_38(2);
ELSE
	BUSLINE(2) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_39)
BEGIN
if (SYNTHESIZED_WIRE_39 = '1') THEN
	BUSLINE(1) <= SYNTHESIZED_WIRE_38(1);
ELSE
	BUSLINE(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_39)
BEGIN
if (SYNTHESIZED_WIRE_39 = '1') THEN
	BUSLINE(0) <= SYNTHESIZED_WIRE_38(0);
ELSE
	BUSLINE(0) <= 'Z';
END IF;
END PROCESS;


b2v_IR : reg16-tri-b-n
PORT MAP(WN => SYNTHESIZED_WIRE_40,
		 RN => SYNTHESIZED_WIRE_41,
		 CLK => SYNTHESIZED_WIRE_62,
		 I => BUSLINE,
		 O => irb);


b2v_MAR : reg16-tri-b-n
PORT MAP(WN => SYNTHESIZED_WIRE_43,
		 RN => SYNTHESIZED_WIRE_44,
		 CLK => SYNTHESIZED_WIRE_62,
		 I => BUSLINE,
		 O => MARB);


PROCESS(SYNTHESIZED_WIRE_62,SYNTHESIZED_WIRE_46)
BEGIN
IF (SYNTHESIZED_WIRE_46 = '0') THEN
	DFF_odff <= '0';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_62)) THEN
	DFF_odff <= halo;
END IF;
END PROCESS;


b2v_PC : reg16-tri-imm-bn
PORT MAP(WN => SYNTHESIZED_WIRE_48,
		 RN => RDPC,
		 CLK => SYNTHESIZED_WIRE_62,
		 D => BUSLINE,
		 Oimm => PC_v,
		 Otri => BUSLINE);


b2v_RAM : ram0
PORT MAP(wren => SYNTHESIZED_WIRE_50,
		 rden => SYNTHESIZED_WIRE_51,
		 inclock => SYNTHESIZED_WIRE_62,
		 address => MARB(7 DOWNTO 0),
		 data => BUSLINE,
		 q => SYNTHESIZED_WIRE_38);


b2v_spA : reg16-tri-imm-bn
PORT MAP(WN => SYNTHESIZED_WIRE_53,
		 RN => SYNTHESIZED_WIRE_54,
		 CLK => SYNTHESIZED_WIRE_62,
		 D => BUSLINE,
		 Oimm => SPAB,
		 Otri => BUSLINE);


b2v_spB : reg16-tri-imm-bn
PORT MAP(WN => SYNTHESIZED_WIRE_56,
		 RN => SYNTHESIZED_WIRE_57,
		 CLK => SYNTHESIZED_WIRE_62,
		 D => BUSLINE,
		 Oimm => SYNTHESIZED_WIRE_32,
		 Otri => BUSLINE);


b2v_spC : reg16-tri-imm-bn
PORT MAP(WN => SYNTHESIZED_WIRE_59,
		 RN => SYNTHESIZED_WIRE_60,
		 CLK => SYNTHESIZED_WIRE_62,
		 D => BUSLINE,
		 Oimm => SYNTHESIZED_WIRE_33,
		 Otri => BUSLINE);

MAR_v(7 DOWNTO 0) <= MARB(7 DOWNTO 0);

END bdf_type;